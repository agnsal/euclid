-- ../../i8051ISS/euclidKeil/Objects/euclid.hex_EOL.hex 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use WORK.I8051_LIB.all;

entity I8051_ROM is
    port(rst      : in  STD_LOGIC;
         clk      : in  STD_LOGIC;
         addr     : in  UNSIGNED (11 downto 0);
         data     : out UNSIGNED (7 downto 0);
         rd       : in  STD_LOGIC);
end I8051_ROM;

architecture BHV of I8051_ROM is

    type ROM_TYPE is array (0 to 2300) of UNSIGNED (7 downto 0);

    constant PROGRAM : ROM_TYPE := (

	"00000010",	-- LJMP   
	"00001000",
	"11101111",
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"00000000",	-- NOP    
	"11000010",	-- CLR_3  
	"11010101",
	"11101100",	-- MOV_1  
	"00110000",	-- JNB    
	"11100111",
	"00001001",
	"10110010",	-- CPL_3  
	"11010101",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10011101",	-- SUBB_1 
	"11111101",	-- MOV_5  
	"11100100",	-- CLR_1  
	"10011100",	-- SUBB_1 
	"11111100",	-- MOV_5  
	"11101110",	-- MOV_1  
	"00110000",	-- JNB    
	"11100111",
	"00010101",
	"10110010",	-- CPL_3  
	"11010101",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10011111",	-- SUBB_1 
	"11111111",	-- MOV_5  
	"11100100",	-- CLR_1  
	"10011110",	-- SUBB_1 
	"11111110",	-- MOV_5  
	"00010010",	-- LCALL  
	"00001000",
	"00110110",
	"11000011",	-- CLR_2  
	"11100100",	-- CLR_1  
	"10011101",	-- SUBB_1 
	"11111101",	-- MOV_5  
	"11100100",	-- CLR_1  
	"10011100",	-- SUBB_1 
	"11111100",	-- MOV_5  
	"10000000",	-- SJMP   
	"00000011",
	"00010010",	-- LCALL  
	"00001000",
	"00110110",
	"00110000",	-- JNB    
	"11010101",
	"00000111",
	"11000011",	-- CLR_2  
	"11100100",	-- CLR_1  
	"10011111",	-- SUBB_1 
	"11111111",	-- MOV_5  
	"11100100",	-- CLR_1  
	"10011110",	-- SUBB_1 
	"11111110",	-- MOV_5  
	"00100010",	-- RET    
	"10111100",	-- CJNE_3 
	"00000000",
	"00001011",
	"10111110",	-- CJNE_3 
	"00000000",
	"00101001",
	"11101111",	-- MOV_1  
	"10001101",	-- MOV_9  
	"11110000",
	"10000100",	-- DIV    
	"11111111",	-- MOV_5  
	"10101101",	-- MOV_6  
	"11110000",
	"00100010",	-- RET    
	"11100100",	-- CLR_1  
	"11001100",	-- XCH_1  
	"11111000",	-- MOV_5  
	"01110101",	-- MOV_12 
	"11110000",
	"00001000",
	"11101111",	-- MOV_1  
	"00101111",	-- ADD_1  
	"11111111",	-- MOV_5  
	"11101110",	-- MOV_1  
	"00110011",	-- RLC    
	"11111110",	-- MOV_5  
	"11101100",	-- MOV_1  
	"00110011",	-- RLC    
	"11111100",	-- MOV_5  
	"11101110",	-- MOV_1  
	"10011101",	-- SUBB_1 
	"11101100",	-- MOV_1  
	"10011000",	-- SUBB_1 
	"01000000",	-- JC     
	"00000101",
	"11111100",	-- MOV_5  
	"11101110",	-- MOV_1  
	"10011101",	-- SUBB_1 
	"11111110",	-- MOV_5  
	"00001111",	-- INC_2  
	"11010101",	-- DJNZ_2 
	"11110000",
	"11101001",
	"11100100",	-- CLR_1  
	"11001110",	-- XCH_1  
	"11111101",	-- MOV_5  
	"00100010",	-- RET    
	"11101101",	-- MOV_1  
	"11111000",	-- MOV_5  
	"11110101",	-- MOV_8  
	"11110000",
	"11101110",	-- MOV_1  
	"10000100",	-- DIV    
	"00100000",	-- JB     
	"11010010",
	"00011100",
	"11111110",	-- MOV_5  
	"10101101",	-- MOV_6  
	"11110000",
	"01110101",	-- MOV_12 
	"11110000",
	"00001000",
	"11101111",	-- MOV_1  
	"00101111",	-- ADD_1  
	"11111111",	-- MOV_5  
	"11101101",	-- MOV_1  
	"00110011",	-- RLC    
	"11111101",	-- MOV_5  
	"01000000",	-- JC     
	"00000111",
	"10011000",	-- SUBB_1 
	"01010000",	-- JNC    
	"00000110",
	"11010101",	-- DJNZ_2 
	"11110000",
	"11110010",
	"00100010",	-- RET    
	"11000011",	-- CLR_2  
	"10011000",	-- SUBB_1 
	"11111101",	-- MOV_5  
	"00001111",	-- INC_2  
	"11010101",	-- DJNZ_2 
	"11110000",
	"11101010",
	"00100010",	-- RET    
	"01111011",	-- MOV_7  
	"01100100",
	"01110101",	-- MOV_12 
	"10000010",
	"00111100",
	"01110101",	-- MOV_12 
	"10000011",
	"00000000",
	"01111111",	-- MOV_7  
	"01100100",
	"01111110",	-- MOV_7  
	"00000000",
	"01111101",	-- MOV_7  
	"00111100",
	"01111100",	-- MOV_7  
	"00000000",
	"00010010",	-- LCALL  
	"00001000",
	"00000000",
	"10001110",	-- MOV_9  
	"00001000",
	"10001111",	-- MOV_9  
	"00001001",
	"01111111",	-- MOV_7  
	"01100100",
	"01111110",	-- MOV_7  
	"00000000",
	"01111101",	-- MOV_7  
	"00111100",
	"01111100",	-- MOV_7  
	"00000000",
	"10000000",	-- SJMP   
	"00101001",
	"11101101",	-- MOV_1  
	"01001100",	-- ORL_1  
	"01100000",	-- JZ     
	"00101010",
	"10001011",	-- MOV_9  
	"10000000",
	"10000101",	-- MOV_10 
	"10000010",
	"10010000",
	"10000101",	-- MOV_10 
	"00001001",
	"10100000",
	"10001101",	-- MOV_9  
	"10110000",
	"10101010",	-- MOV_6  
	"10000011",
	"10101011",	-- MOV_6  
	"10000010",
	"10001100",	-- MOV_9  
	"10000011",
	"10001101",	-- MOV_9  
	"10000010",
	"10101111",	-- MOV_6  
	"00000011",
	"10101110",	-- MOV_6  
	"00000010",
	"00010010",	-- LCALL  
	"00001000",
	"00000000",
	"10001110",	-- MOV_9  
	"00001000",
	"10001111",	-- MOV_9  
	"00001001",
	"10101111",	-- MOV_6  
	"00000011",
	"10101110",	-- MOV_6  
	"00000010",
	"10101101",	-- MOV_6  
	"10000010",
	"10101100",	-- MOV_6  
	"10000011",
	"00010010",	-- LCALL  
	"00001000",
	"00000000",
	"10000000",	-- SJMP   
	"11010010",
	"10001011",	-- MOV_9  
	"10000000",
	"10000101",	-- MOV_10 
	"10000010",
	"10010000",
	"10000101",	-- MOV_10 
	"00001001",
	"10100000",
	"10001101",	-- MOV_9  
	"10110000",
	"11100100",	-- CLR_1  
	"11110101",	-- MOV_8  
	"10000000",
	"11110101",	-- MOV_8  
	"10010000",
	"11110101",	-- MOV_8  
	"10100000",
	"11110101",	-- MOV_8  
	"10110000",
	"10000000",	-- SJMP   
	"11111110",
	"01111000",	-- MOV_7  
	"01111111",
	"11100100",	-- CLR_1  
	"11110110",	-- MOV_13 
	"11011000",	-- DJNZ_1 
	"11111101",
	"01110101",	-- MOV_12 
	"10000001",
	"00001001",
	"00000010",	-- LJMP   
	"00001000",
	"10001011",
	"00000000",	-- NOP    
	"00000000");	-- NOP    
begin

    process(rst, clk)
    begin
        if( rst = '1' ) then

            data <= CD_8;
        elsif( clk'event and clk = '1' ) then

            if( rd = '1' ) then

                data <= PROGRAM(conv_integer(addr));
            else

                data <= CD_8;
            end if;
        end if;
    end process;
end BHV;