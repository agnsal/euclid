-- ../../i8051ISS/euclidSDCC/euclid.hex_EOL.hex 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use WORK.I8051_LIB.all;

entity I8051_ROM is
    port(rst      : in  STD_LOGIC;
         clk      : in  STD_LOGIC;
         addr     : in  UNSIGNED (11 downto 0);
         data     : out UNSIGNED (7 downto 0);
         rd       : in  STD_LOGIC);
end I8051_ROM;

architecture BHV of I8051_ROM is

    type ROM_TYPE is array (0 to 467) of UNSIGNED (7 downto 0);

    constant PROGRAM : ROM_TYPE := (

	"00000010",	-- LJMP   
	"00000000",
	"00000110",
	"00000010",	-- LJMP   
	"00000000",
	"01100010",
	"01110101",	-- MOV_12 
	"10000001",
	"00001001",
	"00010010",	-- LCALL  
	"00000001",
	"11010000",
	"11100101",	-- MOV_2  
	"10000010",
	"01100000",	-- JZ     
	"00000011",
	"00000010",	-- LJMP   
	"00000000",
	"00000011",
	"01111001",	-- MOV_7  
	"00000000",
	"11101001",	-- MOV_1  
	"01000100",	-- ORL_4  
	"00000000",
	"01100000",	-- JZ     
	"00011011",
	"01111010",	-- MOV_7  
	"00000000",
	"10010000",	-- MOV_18 
	"00000001",
	"11010100",
	"01111000",	-- MOV_7  
	"00000001",
	"01110101",	-- MOV_12 
	"10100000",
	"00000000",
	"11100100",	-- CLR_1  
	"10010011",	-- MOVC_1 
	"11110010",	-- MOVX_3 
	"10100011",	-- INC_5  
	"00001000",	-- INC_2  
	"10111000",	-- CJNE_3 
	"00000000",
	"00000010",
	"00000101",	-- INC_3  
	"10100000",
	"11011001",	-- DJNZ_1 
	"11110100",
	"11011010",	-- DJNZ_1 
	"11110010",
	"01110101",	-- MOV_12 
	"10100000",
	"11111111",
	"11100100",	-- CLR_1  
	"01111000",	-- MOV_7  
	"11111111",
	"11110110",	-- MOV_13 
	"11011000",	-- DJNZ_1 
	"11111101",
	"01111000",	-- MOV_7  
	"00000000",
	"11101000",	-- MOV_1  
	"01000100",	-- ORL_4  
	"00000000",
	"01100000",	-- JZ     
	"00001010",
	"01111001",	-- MOV_7  
	"00000001",
	"01110101",	-- MOV_12 
	"10100000",
	"00000000",
	"11100100",	-- CLR_1  
	"11110011",	-- MOVX_3 
	"00001001",	-- INC_2  
	"11011000",	-- DJNZ_1 
	"11111100",
	"01111000",	-- MOV_7  
	"00000000",
	"11101000",	-- MOV_1  
	"01000100",	-- ORL_4  
	"00000000",
	"01100000",	-- JZ     
	"00001100",
	"01111001",	-- MOV_7  
	"00000000",
	"10010000",	-- MOV_18 
	"00000000",
	"00000001",
	"11100100",	-- CLR_1  
	"11110000",	-- MOVX_4 
	"10100011",	-- INC_5  
	"11011000",	-- DJNZ_1 
	"11111100",
	"11011001",	-- DJNZ_1 
	"11111010",
	"00000010",	-- LJMP   
	"00000000",
	"00000011",
	"01111110",	-- MOV_7  
	"01100100",
	"01111111",	-- MOV_7  
	"00000000",
	"01111100",	-- MOV_7  
	"00111100",
	"01111101",	-- MOV_7  
	"00000000",
	"01111010",	-- MOV_7  
	"00000001",
	"01111011",	-- MOV_7  
	"00000000",
	"01111000",	-- MOV_7  
	"00101000",
	"01111001",	-- MOV_7  
	"00000000",
	"11101000",	-- MOV_1  
	"01001001",	-- ORL_1  
	"01100000",	-- JZ     
	"01100000",
	"10001110",	-- MOV_9  
	"10000000",
	"10001100",	-- MOV_9  
	"10010000",
	"10001010",	-- MOV_9  
	"10100000",
	"10001000",	-- MOV_9  
	"10110000",
	"10001100",	-- MOV_9  
	"00000110",
	"10001101",	-- MOV_9  
	"00000111",
	"10001000",	-- MOV_9  
	"00000100",
	"10001001",	-- MOV_9  
	"00000101",
	"10001000",	-- MOV_9  
	"00001000",
	"10001001",	-- MOV_9  
	"00001001",
	"10001110",	-- MOV_9  
	"10000010",
	"10001111",	-- MOV_9  
	"10000011",
	"11000000",	-- PUSH   
	"00000111",
	"11000000",	-- PUSH   
	"00000110",
	"11000000",	-- PUSH   
	"00000101",
	"11000000",	-- PUSH   
	"00000100",
	"11000000",	-- PUSH   
	"00000001",
	"11000000",	-- PUSH   
	"00000000",
	"00010010",	-- LCALL  
	"00000001",
	"10011000",
	"10101010",	-- MOV_6  
	"10000010",
	"10101011",	-- MOV_6  
	"10000011",
	"11010000",	-- POP    
	"00000000",
	"11010000",	-- POP    
	"00000001",
	"11010000",	-- POP    
	"00000100",
	"11010000",	-- POP    
	"00000101",
	"11010000",	-- POP    
	"00000110",
	"11010000",	-- POP    
	"00000111",
	"10001000",	-- MOV_9  
	"00001000",
	"10001001",	-- MOV_9  
	"00001001",
	"10001110",	-- MOV_9  
	"10000010",
	"10001111",	-- MOV_9  
	"10000011",
	"11000000",	-- PUSH   
	"00000111",
	"11000000",	-- PUSH   
	"00000110",
	"11000000",	-- PUSH   
	"00000101",
	"11000000",	-- PUSH   
	"00000100",
	"11000000",	-- PUSH   
	"00000011",
	"11000000",	-- PUSH   
	"00000010",
	"00010010",	-- LCALL  
	"00000001",
	"01100010",
	"10101000",	-- MOV_6  
	"10000010",
	"10101001",	-- MOV_6  
	"10000011",
	"11010000",	-- POP    
	"00000010",
	"11010000",	-- POP    
	"00000011",
	"11010000",	-- POP    
	"00000100",
	"11010000",	-- POP    
	"00000101",
	"11010000",	-- POP    
	"00000110",
	"11010000",	-- POP    
	"00000111",
	"10000000",	-- SJMP   
	"10011100",
	"10001110",	-- MOV_9  
	"10000000",
	"10001100",	-- MOV_9  
	"10010000",
	"10001010",	-- MOV_9  
	"10100000",
	"10001000",	-- MOV_9  
	"10110000",
	"01110101",	-- MOV_12 
	"10000000",
	"00000000",
	"01110101",	-- MOV_12 
	"10010000",
	"00000000",
	"01110101",	-- MOV_12 
	"10100000",
	"00000000",
	"01110101",	-- MOV_12 
	"10110000",
	"00000000",
	"10000000",	-- SJMP   
	"11111110",
	"11100101",	-- MOV_2  
	"00001000",
	"01000101",	-- ORL_2  
	"00001001",
	"01100000",	-- JZ     
	"01000110",
	"01111010",	-- MOV_7  
	"00000001",
	"11100101",	-- MOV_2  
	"00001000",
	"00100101",	-- ADD_2  
	"11100000",
	"11110101",	-- MOV_8  
	"00001000",
	"11100101",	-- MOV_2  
	"00001001",
	"00110011",	-- RLC    
	"01000000",	-- JC     
	"00010010",
	"11110101",	-- MOV_8  
	"00001001",
	"11100101",	-- MOV_2  
	"10000010",
	"10010101",	-- SUBB_2 
	"00001000",
	"11100101",	-- MOV_2  
	"10000011",
	"10010101",	-- SUBB_2 
	"00001001",
	"01000000",	-- JC     
	"00000011",
	"00001010",	-- INC_2  
	"10000000",	-- SJMP   
	"11100110",
	"11000011",	-- CLR_2  
	"11100101",	-- MOV_2  
	"00001001",
	"00010011",	-- RRC    
	"11110101",	-- MOV_8  
	"00001001",
	"11100101",	-- MOV_2  
	"00001000",
	"00010011",	-- RRC    
	"11110101",	-- MOV_8  
	"00001000",
	"11000011",	-- CLR_2  
	"11100101",	-- MOV_2  
	"10000010",
	"10010101",	-- SUBB_2 
	"00001000",
	"11110101",	-- MOV_8  
	"11110000",
	"11100101",	-- MOV_2  
	"10000011",
	"10010101",	-- SUBB_2 
	"00001001",
	"01000000",	-- JC     
	"00000101",
	"11110101",	-- MOV_8  
	"10000011",
	"10000101",	-- MOV_10 
	"11110000",
	"10000010",
	"11000011",	-- CLR_2  
	"11100101",	-- MOV_2  
	"00001001",
	"00010011",	-- RRC    
	"11110101",	-- MOV_8  
	"00001001",
	"11100101",	-- MOV_2  
	"00001000",
	"00010011",	-- RRC    
	"11110101",	-- MOV_8  
	"00001000",
	"11011010",	-- DJNZ_1 
	"11100001",
	"00100010",	-- RET    
	"01111010",	-- MOV_7  
	"00010000",
	"11100100",	-- CLR_1  
	"11111011",	-- MOV_5  
	"11111100",	-- MOV_5  
	"11100101",	-- MOV_2  
	"10000010",
	"00100101",	-- ADD_2  
	"11100000",
	"11110101",	-- MOV_8  
	"10000010",
	"11100101",	-- MOV_2  
	"10000011",
	"00110011",	-- RLC    
	"11110101",	-- MOV_8  
	"10000011",
	"11101011",	-- MOV_1  
	"00110011",	-- RLC    
	"11111011",	-- MOV_5  
	"11101100",	-- MOV_1  
	"00110011",	-- RLC    
	"11111100",	-- MOV_5  
	"11101011",	-- MOV_1  
	"10010101",	-- SUBB_2 
	"00001000",
	"11110101",	-- MOV_8  
	"11110000",
	"11101100",	-- MOV_1  
	"10010101",	-- SUBB_2 
	"00001001",
	"01000000",	-- JC     
	"00000110",
	"11111100",	-- MOV_5  
	"10101011",	-- MOV_6  
	"11110000",
	"01000011",	-- ORL_6  
	"10000010",
	"00000001",
	"11011010",	-- DJNZ_1 
	"11011101",
	"00100010",	-- RET    
	"11000010",	-- CLR_3  
	"11010101",
	"11100101",	-- MOV_2  
	"10000011",
	"00110000",	-- JNB    
	"11100111",
	"00001101",
	"11010010",	-- SETB_2 
	"11010101",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10010101",	-- SUBB_2 
	"10000010",
	"11110101",	-- MOV_8  
	"10000010",
	"11100100",	-- CLR_1  
	"10010101",	-- SUBB_2 
	"10000011",
	"11110101",	-- MOV_8  
	"10000011",
	"11100101",	-- MOV_2  
	"00001001",
	"00110000",	-- JNB    
	"11100111",
	"00001011",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10010101",	-- SUBB_2 
	"00001000",
	"11110101",	-- MOV_8  
	"00001000",
	"11100100",	-- CLR_1  
	"10010101",	-- SUBB_2 
	"00001001",
	"11110101",	-- MOV_8  
	"00001001",
	"00010010",	-- LCALL  
	"00000000",
	"11101100",
	"00110000",	-- JNB    
	"11010101",
	"00001011",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10010101",	-- SUBB_2 
	"10000010",
	"11110101",	-- MOV_8  
	"10000010",
	"11100100",	-- CLR_1  
	"10010101",	-- SUBB_2 
	"10000011",
	"11110101",	-- MOV_8  
	"10000011",
	"00100010",	-- RET    
	"11000010",	-- CLR_3  
	"11010101",
	"11100101",	-- MOV_2  
	"10000011",
	"00110000",	-- JNB    
	"11100111",
	"00001101",
	"11010010",	-- SETB_2 
	"11010101",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10010101",	-- SUBB_2 
	"10000010",
	"11110101",	-- MOV_8  
	"10000010",
	"11100100",	-- CLR_1  
	"10010101",	-- SUBB_2 
	"10000011",
	"11110101",	-- MOV_8  
	"10000011",
	"11100101",	-- MOV_2  
	"00001001",
	"00110000",	-- JNB    
	"11100111",
	"00001101",
	"10110010",	-- CPL_3  
	"11010101",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10010101",	-- SUBB_2 
	"00001000",
	"11110101",	-- MOV_8  
	"00001000",
	"11100100",	-- CLR_1  
	"10010101",	-- SUBB_2 
	"00001001",
	"11110101",	-- MOV_8  
	"00001001",
	"00010010",	-- LCALL  
	"00000001",
	"00111001",
	"00110000",	-- JNB    
	"11010101",
	"00001011",
	"11100100",	-- CLR_1  
	"11000011",	-- CLR_2  
	"10010101",	-- SUBB_2 
	"10000010",
	"11110101",	-- MOV_8  
	"10000010",
	"11100100",	-- CLR_1  
	"10010101",	-- SUBB_2 
	"10000011",
	"11110101",	-- MOV_8  
	"10000011",
	"00100010",	-- RET    
	"01110101",	-- MOV_12 
	"10000010",
	"00000000",
	"00100010");	-- RET    
begin

    process(rst, clk)
    begin
        if( rst = '1' ) then

            data <= CD_8;
        elsif( clk'event and clk = '1' ) then

            if( rd = '1' ) then

                data <= PROGRAM(conv_integer(addr));
            else

                data <= CD_8;
            end if;
        end if;
    end process;
end BHV;